module menorigual_640(x,menor);
	input [9:0]x;
	output menor;
	
	//COMPARAR BIT A BIT
	igual_1bit EQ9(.a(x[9]), .b(1'b1), .saida(igual9));
	igual_1bit EQ8(.a(x[8]), .b(1'b0), .saida(igual8));
	igual_1bit EQ7(.a(x[7]), .b(1'b1), .saida(igual7));
	igual_1bit EQ6(.a(x[6]), .b(1'b0), .saida(igual6));
	igual_1bit EQ5(.a(x[5]), .b(1'b0), .saida(igual5));
	igual_1bit EQ4(.a(x[4]), .b(1'b0), .saida(igual4));
	igual_1bit EQ3(.a(x[3]), .b(1'b0), .saida(igual3));
	igual_1bit EQ2(.a(x[2]), .b(1'b0), .saida(igual2));
	igual_1bit EQ1(.a(x[1]), .b(1'b0), .saida(igual1));
	igual_1bit EQ0(.a(x[0]), .b(1'b0), .saida(igual0));

	// COMPARANDO MENORES
	menor_1bit M9(.a(x[9]), .b(1'b1), .saida(menor9));
	menor_1bit M8(.a(x[8]), .b(1'b0), .saida(menor8));
	menor_1bit M7(.a(x[7]), .b(1'b1), .saida(menor7));
	menor_1bit M6(.a(x[6]), .b(1'b0), .saida(menor6));
	menor_1bit M5(.a(x[5]), .b(1'b0), .saida(menor5));
	menor_1bit M4(.a(x[4]), .b(1'b0), .saida(menor4));
	menor_1bit M3(.a(x[3]), .b(1'b0), .saida(menor3));
	menor_1bit M2(.a(x[2]), .b(1'b0), .saida(menor2));
	menor_1bit M1(.a(x[1]), .b(1'b0), .saida(menor1));
	menor_1bit M0(.a(x[0]), .b(1'b0), .saida(menor0));
	
	// DEFINIR QUANDO E MENOR POR NIVEL
	and (nivel8,igual9,menor8);
	and(nivel7)
	or (menor,menor9,nivel8)

endmodule



module TOP_MODULE (A,B,C,D,E, Disp1, Disp2, Disp3, LED);
    input A,B,C,D,E;
    output [6:0]Disp1, Disp2, Disp3, LED;
    wire C1;  // Carry entre os dois somadores de 1 bit

    // Instanciando o primeiro somador completo de 1 bit (bit menos significativo)
    HexaMaiSig DISPLAY02 (
        .A(A),
        .B(B),
        .C(C),
        .D(D),
		  .E(E),
        .segA(Disp2[0]),
		  .segB(Disp2[1]),
		  .segC(Disp2[2]),
		  .segD(Disp2[3]),
		  .segE(Disp2[4]),
		  .segF(Disp2[5]),
		  .segG(Disp2[6])
    );

    // Instanciando o segundo somador completo de 1 bit (bit mais significativo)
     HexaMenoSig DISPLAY01 (
        .A(A),
        .B(B),
        .C(C),
        .D(D),
		  .E(E),
        .segA(Disp1[0]),
		  .segB(Disp1[1]),
		  .segC(Disp1[2]),
		  .segD(Disp1[3]),
		  .segE(Disp1[4]),
		  .segF(Disp1[5]),
		  .segG(Disp1[6])
    );
	 
	 caractere DISPLAY03 (
			.A(A),
			.B(B),
			.C(C),
			.D(D),
			.E(E),
			.a(Disp3[0]),
			.b(Disp3[1]),
			.c(Disp3[2]),
			.d(Disp3[3]),
			.e(Disp3[4]),
			.f(Disp3[5]),
			.g(Disp3[6])
	);
	
	binario LEDS (
			.A(A),
			.B(B),
			.C(C),
			.D(D),
			.E(E),
			.S6(LED[6]),
			.S5(LED[5]),
			.S4(LED[4]),
			.S3(LED[3]),
			.S2(LED[2]),
			.S1(LED[1]),
			.S0(LED[0]) 
	);
			

endmodule