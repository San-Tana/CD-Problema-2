module igual_1bit( input a, input b, output saida);
	xnor(saida,a,b);
endmodule