module soma_10bit(input [9:0] a, input [9:0] b, output [9:0] s);
    wire c1, c2, c3, c4, c5, c6, c7, c8, c9;

    full_adder f0(a[0], b[0], 1'b0,  s[0], c1);
    full_adder f1(a[1], b[1], c1,    s[1], c2);
    full_adder f2(a[2], b[2], c2,    s[2], c3);
    full_adder f3(a[3], b[3], c3,    s[3], c4);
    full_adder f4(a[4], b[4], c4,    s[4], c5);
	 
	 full_adder f5(a[5], b[5], c5,    s[5], c6);
	 full_adder f6(a[6], b[6], c6,    s[6], c7);
	 full_adder f7(a[7], b[7], c7,    s[7], c8);
	 full_adder f8(a[8], b[8], c8,    s[8], c9);
	 full_adder f9(a[9], b[9], c9,    s[9], /*ignora carry final*/);

endmodule

module full_adder(input a, input b, input cin, output s, output cout);
    wire s1, c1, c2, c3;
    xor(s1, a, b);
    xor(s, s1, cin);
    and(c1, a, b);
    and(c2, a, cin);
    and(c3, b, cin);
    or(cout, c1, c2, c3);
endmodule
